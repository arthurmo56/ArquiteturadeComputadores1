/*

Guia_0402.v
Aluno- Arthur Martinho Medeiros Oliveira	
Matricula- 813168

*/
module Simplified_e(output f, input x, y);
assign f = ~y & ~x;
endmodule
